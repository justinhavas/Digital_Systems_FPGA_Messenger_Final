module product_register(clk,we,d,res,q);
input clk, we, res;
	input [63:0] d;
	output [63:0] q;
	wire en;
	
	and and1(en,clk,we);
	dffe_ref dff0(q[0],d[0],clk,en,res);
	dffe_ref dff1(q[1],d[1],clk,en,res);
	dffe_ref dff2(q[2],d[2],clk,en,res);
	dffe_ref dff3(q[3],d[3],clk,en,res);
	dffe_ref dff4(q[4],d[4],clk,en,res);
	dffe_ref dff5(q[5],d[5],clk,en,res);
	dffe_ref dff6(q[6],d[6],clk,en,res);
	dffe_ref dff7(q[7],d[7],clk,en,res);
	dffe_ref dff8(q[8],d[8],clk,en,res);
	dffe_ref dff9(q[9],d[9],clk,en,res);
	dffe_ref dff10(q[10],d[10],clk,en,res);
	dffe_ref dff11(q[11],d[11],clk,en,res);
	dffe_ref dff12(q[12],d[12],clk,en,res);
	dffe_ref dff13(q[13],d[13],clk,en,res);
	dffe_ref dff14(q[14],d[14],clk,en,res);
	dffe_ref dff15(q[15],d[15],clk,en,res);
	dffe_ref dff16(q[16],d[16],clk,en,res);
	dffe_ref dff17(q[17],d[17],clk,en,res);
	dffe_ref dff18(q[18],d[18],clk,en,res);
	dffe_ref dff19(q[19],d[19],clk,en,res);
	dffe_ref dff20(q[20],d[20],clk,en,res);
	dffe_ref dff21(q[21],d[21],clk,en,res);
	dffe_ref dff22(q[22],d[22],clk,en,res);
	dffe_ref dff23(q[23],d[23],clk,en,res);
	dffe_ref dff24(q[24],d[24],clk,en,res);
	dffe_ref dff25(q[25],d[25],clk,en,res);
	dffe_ref dff26(q[26],d[26],clk,en,res);
	dffe_ref dff27(q[27],d[27],clk,en,res);
	dffe_ref dff28(q[28],d[28],clk,en,res);
	dffe_ref dff29(q[29],d[29],clk,en,res);
	dffe_ref dff30(q[30],d[30],clk,en,res);
	dffe_ref dff31(q[31],d[31],clk,en,res);
	dffe_ref dff32(q[32],d[32],clk,en,res);
	dffe_ref dff33(q[33],d[33],clk,en,res);
	dffe_ref dff34(q[34],d[34],clk,en,res);
	dffe_ref dff35(q[35],d[35],clk,en,res);
	dffe_ref dff36(q[36],d[36],clk,en,res);
	dffe_ref dff37(q[37],d[37],clk,en,res);
	dffe_ref dff38(q[38],d[38],clk,en,res);
	dffe_ref dff39(q[39],d[39],clk,en,res);
	dffe_ref dff40(q[40],d[40],clk,en,res);
	dffe_ref dff41(q[41],d[41],clk,en,res);
	dffe_ref dff42(q[42],d[42],clk,en,res);
	dffe_ref dff43(q[43],d[43],clk,en,res);
	dffe_ref dff44(q[44],d[44],clk,en,res);
	dffe_ref dff45(q[45],d[45],clk,en,res);
	dffe_ref dff46(q[46],d[46],clk,en,res);
	dffe_ref dff47(q[47],d[47],clk,en,res);
	dffe_ref dff48(q[48],d[48],clk,en,res);
	dffe_ref dff49(q[49],d[49],clk,en,res);
	dffe_ref dff50(q[50],d[50],clk,en,res);
	dffe_ref dff51(q[51],d[51],clk,en,res);
	dffe_ref dff52(q[52],d[52],clk,en,res);
	dffe_ref dff53(q[53],d[53],clk,en,res);
	dffe_ref dff54(q[54],d[54],clk,en,res);
	dffe_ref dff55(q[55],d[55],clk,en,res);
	dffe_ref dff56(q[56],d[56],clk,en,res);
	dffe_ref dff57(q[57],d[57],clk,en,res);
	dffe_ref dff58(q[58],d[58],clk,en,res);
	dffe_ref dff59(q[59],d[59],clk,en,res);
	dffe_ref dff60(q[60],d[60],clk,en,res);
	dffe_ref dff61(q[61],d[61],clk,en,res);
	dffe_ref dff62(q[62],d[62],clk,en,res);
	dffe_ref dff63(q[63],d[63],clk,en,res);
endmodule