module not_bitwise(in1,out);
	input [31:0] in1;
	output [31:0] out;
	
	not not0(out[0],in1[0]);
	not not1(out[1],in1[1]);
	not not2(out[2],in1[2]);
	not not3(out[3],in1[3]);
	not not4(out[4],in1[4]);
	not not5(out[5],in1[5]);
	not not6(out[6],in1[6]);
	not not7(out[7],in1[7]);
	not not8(out[8],in1[8]);
	not not9(out[9],in1[9]);
	not not10(out[10],in1[10]);
	not not11(out[11],in1[11]);
	not not12(out[12],in1[12]);
	not not13(out[13],in1[13]);
	not not14(out[14],in1[14]);
	not not15(out[15],in1[15]);
	not not16(out[16],in1[16]);
	not not17(out[17],in1[17]);
	not not18(out[18],in1[18]);
	not not19(out[19],in1[19]);
	not not20(out[20],in1[20]);
	not not21(out[21],in1[21]);
	not not22(out[22],in1[22]);
	not not23(out[23],in1[23]);
	not not24(out[24],in1[24]);
	not not25(out[25],in1[25]);
	not not26(out[26],in1[26]);
	not not27(out[27],in1[27]);
	not not28(out[28],in1[28]);
	not not29(out[29],in1[29]);
	not not30(out[30],in1[30]);
	not not31(out[31],in1[31]);
endmodule